--------------------------------------------------------------------------------
-- r-VEX | Instruction ROM
--------------------------------------------------------------------------------
-- 
-- This file was assembled by r-ASM, the r-VEX assembler/
-- instruction ROM generator.
-- 
--     source file: ../../demos/fibonacci.s
--     r-ASM flags: ./rasm ../../demos/fibonacci.s
--     date & time: Jul 19, 2008 @ 17:01:38
-- 
-- r-VEX & r-ASM are
-- Copyright (c) 2008, Thijs van As <t.vanas@gmail.com>
-- 
-- Computer Engineering Laboratory
-- Delft University of Technology
-- Delft, The Netherlands
-- 
-- http://r-vex.googlecode.com
-- 
-- r-VEX is free hardware: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
-- 
--------------------------------------------------------------------------------
-- i_mem.vhd (generated by r-ASM)
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity i_mem is
	port ( reset   : in std_logic;                        -- system reset
	       address : in std_logic_vector(7 downto 0);     -- address of instruction to be read

	       instr   : out std_logic_vector(127 downto 0)); -- instruction (4 syllables)
end entity i_mem;


architecture behavioural of i_mem is
begin
	memory : process(address, reset)
	begin
		if (reset = '1') then
			instr <= x"00000000000000000000000000000000";
		else
			case address is
				when x"00"  => instr <= "10000011000111100000000000000110"& -- add $r0.15 = $r0.0, 1
				                        "10110000000000100000000000000000"& -- mov $r0.1 = $r0.0
				                        "10000011000101000000000010110000"& -- add $r0.10 = $r0.0, 44
				                        "10000011000001000000000000000101"; -- add $r0.2 = $r0.0, 1
				                                                            -- LABEL_BEGIN:
				when x"01"  => instr <= "10000010000001000000100001000010"& -- add $r0.2 = $r0.1, $r0.2
				                        "10000010000001100000000001000000"& -- add $r0.3 = $r0.0, $r0.2
				                        "10110010000000000100100101000000"& -- cmpeq $b0.0 = $r0.9, $r0.10
				                        "01001010100000000000000001100001"; -- br $b0.0, LABEL_END
				when x"02"  => instr <= "10000011000100100100100000000110"& -- add $r0.9 = $r0.9, 1
				                        "10000010000000100000000001100000"& -- add $r0.1 = $r0.0, $r0.3
				                        "00000000000000000000000000000000"& -- nop
				                        "01000010100000000000000000100001"; -- goto LABEL_BEGIN
				                                                            -- LABEL_END:
				when x"03"  => instr <= "00101100000000100111100000000010"& -- stw 0x0[$r0.15] = $r0.1
				                        "10110000000100100000000000000000"& -- mov $r0.9 = $r0.0
				                        "00000000000000000000000000000000"& -- nop
				                        "00000000000000000000000000000001"; -- nop
				when others => instr <= "00000000000000000000000000000010"& -- nop
				                        "00000000000000000000000000000000"& -- nop
				                        "00000000000000000000000000000000"& -- nop
				                        "00111110000000000000000000000001"; -- stop
			end case;
		end if;
	end process memory;
end architecture behavioural;

